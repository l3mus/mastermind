bit_12_counter_inst : bit_12_counter PORT MAP (
		clock	 => clock_sig,
		cnt_en	 => cnt_en_sig,
		q	 => q_sig
	);
